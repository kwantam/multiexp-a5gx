localparam CMD_BEGINRAMMULT = 3'b001;
localparam CMD_BEGINMULT    = 3'b010;
localparam CMD_BEGINSQUARE  = 3'b011;
localparam CMD_PRELOAD      = 3'b100;
localparam CMD_STORE        = 3'b101;
localparam CMD_RESETRESULT  = 3'b110;
localparam CMD_INVALID      = 3'b111;
